
module RCA_16_bit(input logic [15:0]a,b,output logic [16:0]s

    );
    logic [14:0]c;
   fa f1(a[0],b[0],1'b0,s[0],c[0]);
   fa f2(a[1],b[1],c[0],s[1],c[1]);
   fa f3(a[2],b[2],c[1],s[2],c[2]);
   fa f4(a[3],b[3],c[2],s[3],c[3]);
   fa f5(a[4],b[4],c[3],s[4],c[4]);
   fa f6(a[5],b[5],c[4],s[5],c[5]);
   fa f7(a[6],b[6],c[5],s[6],c[6]);
   fa f8(a[7],b[7],c[6],s[7],c[7]);
   fa f9(a[8],b[8],c[7],s[8],c[8]);
   fa f10(a[9],b[9],c[8],s[9],c[9]);
   fa f11(a[10],b[10],c[9],s[10],c[10]);
   fa f12(a[11],b[11],c[10],s[11],c[11]);
   fa f13(a[12],b[12],c[11],s[12],c[12]);
   fa f14(a[13],b[13],c[12],s[13],c[13]);
   fa f15(a[14],b[14],c[13],s[14],c[14]);
   fa f16(a[15],b[15],c[14],s[15],s[16]);
   
endmodule
