
module broun_multi(input logic [7:0]a,b,output logic [15:0]y

    );
    logic[56:1]s,c;
    logic p[7:0][7:0];
    always_comb
    begin
    for(int i=0;i<=7;i++) 
      for(int j=0;j<=7;j++)
         p[j][i]<=a[j]&b[i];
    end
    //first line
    fa f1(p[1][0],p[0][1],1'b0,s[1],c[1]);
    fa f2(p[2][0],p[1][1],c[1],s[2],c[2]);
    fa f3(p[3][0],p[2][1],c[2],s[3],c[3]);
    fa f4(p[4][0],p[3][1],c[3],s[4],c[4]);
    fa f5(p[5][0],p[4][1],c[4],s[5],c[5]);
    fa f6(p[6][0],p[5][1],c[5],s[6],c[6]);
    fa f7(p[7][0],p[6][1],c[6],s[7],c[7]);
    fa f8(1'b0,p[7][1],c[7],s[8],c[8]);
    //second line
    fa f9(s[2],p[0][2],1'b0,s[9],c[9]);
    fa f10(s[3],p[1][2],c[9],s[10],c[10]);
    fa f11(s[4],p[2][2],c[10],s[11],c[11]);
    fa f12(s[5],p[3][2],c[11],s[12],c[12]);
    fa f13(s[6],p[4][2],c[12],s[13],c[13]);
    fa f14(s[7],p[5][2],c[13],s[14],c[14]);
    fa f15(s[8],p[6][2],c[14],s[15],c[15]);
    fa f16(c[8],p[7][2],c[15],s[16],c[16]);
    //third line
    fa f17(s[10],p[0][3],1'b0,s[17],c[17]);
    fa f18(s[11],p[1][3],c[17],s[18],c[18]);
    fa f19(s[12],p[2][3],c[18],s[19],c[19]);
    fa f20(s[13],p[3][3],c[19],s[20],c[20]);
    fa f21(s[14],p[4][3],c[20],s[21],c[21]);
    fa f22(s[15],p[5][3],c[21],s[22],c[22]);
    fa f23(s[16],p[6][3],c[22],s[23],c[23]);
    fa f24(c[16],p[7][3],c[23],s[24],c[24]);
    //fourth line
    fa f25(s[18],p[0][4],1'b0,s[25],c[25]);
    fa f26(s[19],p[1][4],c[25],s[26],c[26]);
    fa f27(s[20],p[2][4],c[26],s[27],c[27]);
    fa f28(s[21],p[3][4],c[27],s[28],c[28]);
    fa f29(s[22],p[4][4],c[28],s[29],c[29]);
    fa f30(s[23],p[5][4],c[29],s[30],c[30]);
    fa f31(s[24],p[6][4],c[30],s[31],c[31]);
    fa f32(c[24],p[7][4],c[31],s[32],c[32]);
    //fifth line 
    fa f33(s[26],p[0][5],1'b0,s[33],c[33]);
    fa f34(s[27],p[1][5],c[33],s[34],c[34]);
    fa f35(s[28],p[2][5],c[34],s[35],c[35]);
    fa f36(s[29],p[3][5],c[35],s[36],c[36]);
    fa f37(s[30],p[4][5],c[36],s[37],c[37]);
    fa f38(s[31],p[5][5],c[37],s[38],c[38]);
    fa f39(s[32],p[6][5],c[38],s[39],c[39]);
    fa f40(c[32],p[7][5],c[39],s[40],c[40]);
    //six line
    fa f41(s[34],p[0][6],1'b0,s[41],c[41]);
    fa f42(s[35],p[1][6],c[41],s[42],c[42]);
    fa f43(s[36],p[2][6],c[42],s[43],c[43]);
    fa f44(s[37],p[3][6],c[43],s[44],c[44]);
    fa f45(s[38],p[4][6],c[44],s[45],c[45]);
    fa f46(s[39],p[5][6],c[45],s[46],c[46]);
    fa f47(s[40],p[6][6],c[46],s[47],c[47]);
    fa f48(c[40],p[7][6],c[47],s[48],c[48]);
    //seventh line
    fa f49(s[42],p[0][7],1'b0,s[49],c[49]);
    fa f50(s[43],p[1][7],c[49],s[50],c[50]);
    fa f51(s[44],p[2][7],c[50],s[51],c[51]);
    fa f52(s[45],p[3][7],c[51],s[52],c[52]);
    fa f53(s[46],p[4][7],c[52],s[53],c[53]);
    fa f54(s[47],p[5][7],c[53],s[54],c[54]);
    fa f55(s[48],p[6][7],c[54],s[55],c[55]);
    fa f56(c[48],p[7][7],c[55],s[56],c[56]);
       
   assign y[0]=p[0][0]; 
   assign y[1]=s[1]; 
   assign y[2]=s[9]; 
   assign y[3]=s[17]; 
   assign y[4]=s[25]; 
   assign y[5]=s[33]; 
   assign y[6]=s[41]; 
   assign y[7]=s[49]; 
   assign y[8]=s[50]; 
   assign y[9]=s[51]; 
   assign y[10]=s[52]; 
   assign y[11]=s[53]; 
   assign y[12]=s[54]; 
   assign y[13]=s[55]; 
   assign y[14]=s[56]; 
   assign y[15]=c[56]; 
      
endmodule
